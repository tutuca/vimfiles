b0VIM 7.3      !�9M� P<  pandres                                 acerina                                 ~pandres/projects/bixti/kioskito/apps/kiosquero/views/base.py                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                utf-8	 3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           [                            h       \              	       ]       �                     =       !                    !       U                    ]       u                    e       �                    1       7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ad  %   �     [       �  �  m    �  �  z  G  �  �  �  L  %    �  �  �  o  H  G    �  �  w  v  N  �
  
  
  �	  �	  �	  �	  o	  n	  P	  '	  &	  �  �  �  �  �    w  M    �  �  �  �  o  O  5    �  �  �  �  �  �  o  X  +  �  �  �  q  P  9    �  �  }  .    �  �  �  �  k  L     �  �  �    P    �  �  �                                                   shop_config.shipping_countries.clear()             shop_config.in_country_only = False             shop_config.store_name = unicode(data['shop_name'])                 kiosko.banner = data['banner']             if data['banner']:                 kiosko.logo = data['logo']             if data['logo']:             kiosko.site.name = unicode(data['shop_name'])             data = config_form.cleaned_data             kiosko.skin = skin                 skin = kiosko.skin             except:                 skin = Skin.objects.get(slug=request.POST['skin'])             try:             # Kiosko         if config_form.is_valid():                          'banner':request.FILES.get('banner', kiosko.banner)})                         {'logo':request.FILES.get('logo', kiosko.logo),         config_form = ConfigForm(request.POST,         rename_files(request.FILES)     if request.method == 'POST':     config_form = None     skins.insert(0, kiosko.skin)     skins = [skin for skin in skins]     skins = skins.exclude(pk=kiosko.skin.pk)     kiosko = Kiosko.objects.get(site = shop_config.site)     shop_config = Config.objects.get_current()     skins = Skin.objects.filter(active=True)     # Shop Config form def design_store(request): @user_passes_test(is_store_admin)      )         }             'out_of_stock': cnt_out_of_stock             'cnt_products': cnt_products,             'products':products,         extra_context = {         'kiosquero/index.html',         request,     return direct_to_template(          cnt_out_of_stock = len(products.filter(items_in_stock__lte=0))     cnt_products = len(products)     products = Product.objects.filter(site=kiosko.site, active=True)     kiosko = Kiosko.objects.get_current()     '''     Main view of the store management front end.      ''' def index(request): @user_passes_test(is_store_admin)  USER_DELETABLES = (Product, Category, FlatPage, Skin)  log = get_logger('kiosquero.views.base') from logger import get_logger  from decorators import is_store_admin  from shipping_payments import reset_payment_shipping, config_live                              AttributesForm, ConfigDomainForm                             ConfigForm, PageForm, ShopExtrasForm, ConfigStoreForm, GoogleSettingsForm, \ from kiosquero.forms import ProductForm, PriceForm, ProductImageForm, CategoryForm, SellerForm, \ from heladera.models import Customer, Seller, Skin, Plan, Rubro, Kiosko, PaymentMethod, GET_CONFIG_CACHE_KEY from heladera.views import response_add  from l10n.models import Country, AdminArea from livesettings import ConfigurationSettings from product.models import Product, Category, Price, ProductImage from satchmo_store.shop.models import Config, Order  from django.core.mail import send_mail from django.core.cache import cache from django.core.urlresolvers import reverse from django.template import RequestContext from django import forms from django.conf import settings from django.db.models import get_model from django.contrib.flatpages.models import FlatPage from django.contrib.sites.models import Site from django.contrib.auth.decorators import login_required, user_passes_test from django.shortcuts import render_to_response, redirect, get_object_or_404 from django.utils.translation import ugettext as _ from django.utils.encoding import smart_unicode from django.utils import simplejson from django.http import HttpResponse, HttpResponseRedirect, Http404 from django.views.generic.create_update import update_object, create_object, delete_object from django.views.generic.list_detail import object_list, object_detail from django.views.generic.simple import direct_to_template import datetime ad  	  �	     1       �  �  �  �  �  �  �  w  X  G       �  �  �  �  �  �  Q    �  �  �  �  X      �  �  x  0  	  �  �  n  m  )      �
  �
  �
  �
  �
  ;
  �	  �	  �	  �	  �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         files[k].name += datetime.datetime.now().strftime("%Y%m%d%H%M%S%f")         files[k].name = files[k].name.encode('ascii', 'ignore').replace(' ', '_')     for k in files.keys(): def rename_files(files):            return JSONResponse({'error': 'Not Ajax or no GET'})     else:             for o in states])         return JSONResponse([{'id': o.id, 'name': smart_unicode(o)}              cache.set(states_key, states, settings.CACHE_TIMEOUT)             states = AdminArea.objects.filter(country=country_id)         if not states:         states = cache.get(states_key)         states_key = "states_for_country_%(id)s" % {'id': country_id, }         country_id = request.GET['country_id']     if request.is_ajax() and request.GET and 'country_id' in request.GET: def states_for_country(request):                  simplejson.dumps(data), mimetype='application/json')         super(JSONResponse, self).__init__(     def __init__(self, data): class JSONResponse(HttpResponse):                         special=('_thanksstore', reverse(thanks_store)))                        template='mostrador/product_form_step.html',                        product_slug=product_slug,     return new_product(request, def new_product_step(request, product_slug=None): @user_passes_test(is_store_admin)      )         }         extra_context={         'kiosquero/thanks_store.html',         request,     return direct_to_template( def thanks_store(request): @user_passes_test(is_store_admin)       )         }             'form':extra_form,             'skins':skins, ad    (     =       �  �  y  ?    �  �  �  �  z  A  @  2  �  �  �  Q  	  �  �  Q  G  )  �  �  a      �
  �
  �
  d
  c
  <
  
  �	  w	  7	  �  �  X  '  &     �  �  b  a  M  +    �  �  �  <  -  �  �  i  )  (  �  �  �  �  /  �  �  Y  "  �  �  |  g  =  �  �  u  ,      �  �  }  |                       ret_path = request.GET.get('return', reverse('manage')) def delete_by_id(request, model, pk=None): @user_passes_test(is_store_admin)                            slug=slug)                          return HttpResponse(json, mimetype        return HttpRe        return HttpResponse(json, mimetype='application/json')         json = simplejson.dump        return HttpResponse(json        return HttpResponse(json, mimetyp        return HttpResponse(json, mimetype='application        return HttpResponse(json, mimetype='applicat        return HttpResponse(json, mimetype='application/json')               return HttpResponse(json, mimetype='application/json')         json = simplejson.dump        return HttpResponse(json, mimetype='application/json')         json = simplejson.dumps(results)             return HttpRes                 return H                 return HttpResponse(json         return HttpResponse(json, mimetype='applicat    #     return HttpResponse(json, mimetype='application/json')    #     json = simplejson.dumps(results)    #         results = {'success':False, 'errors':_('The category already exists.')}    #         cat = Category.objects.get(site=kiosko.site, name=name)    #     else:    #         results = {'success':False, 'errors':_('The name of the category is required')}    #     if not name:    #     name = request.GET.get(u'category_name', None)    # elif request.is_ajax(): def delete(request, model, slug=None): @user_passes_test(is_store_admin) ## delete Views                                     'form.html')     return direct_to_template(request,     #FIXME: Try to figure out how to return a formclass based of it's name def render_form(request, form_class):                                                })                                               'image_form':image_form,                                               'attributes_form':attributes_form,                                               'price_form':price_form,                                               'errors': errors,                                               'shop_config':kiosko.get_config(),                                extra_context={'product_form':product_form,                                template,     return direct_to_template(request,              image_form = ProductImageForm()             attributes_form = AttributesForm()             price_form = PriceForm()             product_form = ProductForm()         else :             image_form = ProductImageForm(instance=product_instance)             attributes_form = AttributesForm(instance=product_instance)             price_form = PriceForm(instance=product_instance)             product_form = ProductForm(instance=product_instance)         if product_instance :     else:                                           instance=product_instance)                                           request.FILES,              image_form = ProductImageForm(request.POST,                                               instance=product_instance)             attributes_form = AttributesForm(request.POST,                                     instance=product_instance)             price_form = PriceForm(request.POST,              errors = [_("Correct the errors below")]         else:                  errors = [_("Correct the errors below")]             else:                 return response_add(request, product, special=special)                  image_form.save()                 attributes_form.save()                 price_form.save()                     image_form and image_form.is_valid():             if price_form.is_valid() and attributes_form.is_valid() and \                                            instance=product) ad  �	  y
     !       �  �  '    �  �  �  y  O  5  �  �  i  '  �  �  �  �  �  I      �  �  �  �  q  (      �
  �
  y
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ret_path = request.GET.get('return', reverse('manage')) def delete_by_id(request, model, pk=None): @user_passes_test(is_store_admin)                            slug=slug)                           template_name='kiosquero/confirm_delete.html',                           ret_path,                           modelm,     return delete_object(request,         raise Http404         # fail security test     except:         obj = get_object_or_404(objs, slug=slug)             objs = modelm.objects.filter(owner=request.user)         except:             objs = modelm.objects.filter(site=kiosko.site)         try:                 kiosko.save()                 kiosko.skin = default_skin             for kiosko in Kiosko.objects.filter(skin__slug=slug):             default_skin = Skin.objects.get(slug=settings.DEFAULT_SKIN)         if request.POST.get('post', False) and modelm == Skin:         # assign default skin for kioskos that use the removing skin             raise Http404         if modelm not in USER_DELETABLES:         modelm = get_model(app_name,model)         app_name,model = model.split('.')         kiosko = Kiosko.objects.get_current()     try:         return redirect(ret_path)         request.user.message_set.create(message=_('Nothing to delete, operation cancelled'))     if request.POST and request.POST.get('post', 'no') == 'no':     ret_path = request.GET.get('return', reverse('manage')) ad  F   �     ]       �  c  A  8  
  �  �  �  q  +  �  �  �  �  �  {  W    �  �  �  �  �  G  B  *      �  �  �  �  s  I  ,  �
  �
  �
  �
  �
  a
  
  
  �	  �	  �	  b	  F	  	  �  �  �  O  A  0  �  �  f  Q  �  �  �  t  @  �  �  2    �  �  �  �  L  B  $  �  �  K  =    	  �  �  �  �  W  E  7  6  5       �  �                                                                            kiosko = Kiosko.objects.get_current() def page(request): @user_passes_test(is_store_admin)               )                 }                     'form':category_form,                 extra_context={                 'kiosquero/category_form.html',                 request,     return direct_to_template(                      category_form = CategoryForm()         else:             results = {'success':False, 'errors':_('The category already exists.')}         elif Category.objects.get(site=kiosko.site, name=name):             category_form = CategoryForm(instance=category_instance)         if category_instance:     else:         return HttpResponse(json, mimetype='application/json')         json = simplejson.dumps(results)                      results = {'success':False, 'errors':'%s' %e}                 except Exception, e:                     }                         'url_delete': reverse('delete', args=['product.Category', category_instance.slug]),                         'url_edit': reverse('edit_category', args=[category_instance.slug]),                         'url': category_instance.get_absolute_url(),                         'id': category_instance.id,                         'name':category_instance.name,                         'success':True,                      results = {                     category_instance = Category.objects.create(site=kiosko.site, name=name)                 try:             except Category.DoesNotExist:                 results = {'success':False, 'errors':_('The category already exists.')}                 cat = Category.objects.get(site=kiosko.site, name=name)             try:         else:             results = {'success':False, 'errors':_('The name of the category is required')}         if not name:         name = request.GET.get(u'category_name', None)     elif request.is_ajax():             return response_add(request, category)             category.save()             category.rubro_set = data['rubros']             data = category_form.cleaned_data             category = category_form.save()         if category_form.is_valid():          category_form = CategoryForm(request.POST, instance=category_instance)     if request.method == 'POST':                  category_instance = get_object_or_404(categories, slug=category_slug)     if category_slug:      categories = Category.objects.filter(site=kiosko.site)      category_instance = None     kiosko = Kiosko.objects.get_current() def new_category(request, category_slug=None): @user_passes_test(is_store_admin)      )         template_name='kiosquero/manage_categories.html',         categories,         request,     return object_list(          categories = Category.objects.filter(site=kiosko.site)     kiosko = Kiosko.objects.get_current() def category(request): @user_passes_test(is_store_admin)                            object_id=pk)                           template_name='kiosquero/confirm_delete.html',                           ret_path,                           modelm,     return delete_object(request,         raise Http404         # fail security test     except:         obj = get_object_or_404(objs, pk=pk)         objs = modelm.objects.filter(sites__id__exact=kiosko.site.id)             raise Http404         if modelm not in USER_DELETABLES:         modelm = get_model(app_name,model)         app_name,model = model.split('.')         kiosko = Kiosko.objects.get_current()     try:         return redirect(ret_path)         request.user.message_set.create(message=_('Nothing to delete, operation cancelled'))     if request.POST and request.POST.get('post', 'no') == 'no': ad     �     e       �  �  �  �  ~  I  C  B     �  �  �  r  q  a  $    �  �  �  �  q  1  '    �  �  �  �  q  6  �  �  �  �  �  �  ^  F  )  �
  �
  �
  c
  b
  @
  
  �	  �	  �	  �	  b	  7	  	  �  �  �  �  s  7    �  �  i  8    �  �  }  |  V    �  �  �  L    �  �  ~  O    �  �  �  �  Z  	  �  �  �  �  �  }  V  2  1      �  �  �                            extra_context={         'mostrador/create_store.html',         request,     return direct_to_template(      log.debug('Rendering template')         extra_form = ShopExtrasForm()      else:                          return redirect('new_product_step')                  cat.save()                 cat.rubro_set.add(rubro)                 cat = Category.objects.create(site=kiosko.site, name=rubro.name)             for rubro in kiosko.rubro.all():             # create cateogries using rubros              cache.delete(GET_CONFIG_CACHE_KEY % {'id': kiosko.id})             store_config.save()             store_config.postal_code = data['zipcode']             store_config.phone = data['phone']             store_config.city = data['city']             store_config.state = data['state'].name             store_config.street1 = data['address']             store_config.store_email = kiosko.owner.email                 store_config.shipping_countries.add(country)             for country in data['incountries']:             store_config.shipping_countries.clear()             store_config.in_country_only = False             store_config = Config.objects.get_current()             # save shipping countries                  raise forms.ValidationError('The seller does not exists')             except Exception, e:                 seller.save()                 seller.postcode = data['zipcode']                 seller.telephone = data['phone']                 seller.city = data['city']                 seller.state = data['state'].name                 seller.country = data['country'].printable_name                 seller.address = data['address']                 seller = Seller.objects.from_kiosko(kiosko)             try:                  raise forms.ValidationError('The kiosko does not exists')             except Exception, e:                 kiosko.save()                 kiosko.logo=data['logo']                 kiosko.rubro=data['rubro']                 kiosko.skin=skin                 kiosko = Kiosko.objects.get_current()             try:                         skin = Skin.objects.get(slug=request.POST['skin'])             data = extra_form.cleaned_data         if extra_form.is_valid():          extra_form = ShopExtrasForm(request.POST, request.FILES)         rename_files(request.FILES)     if request.method == 'POST':     #items = Category.objects.filter(name__icontains=q)[:limit]     log.debug('skin loaded')     user = request.user     skins = Skin.objects.filter(active=True)     log.info('Entering to step two view') def create_store(request): @user_passes_test(is_store_admin)                                  extra_context={'form':page_form,})                                'kiosquero/page_form.html',     return direct_to_template(request,                      page_form = PageForm()         else :             page_form = PageForm(instance=page_instance)         if page_instance :     else:             return response_add(request, page, slug_or_id='pk')             page = page_form.save()         if page_form.is_valid():          page_form = PageForm(request.POST, instance=page_instance)     if request.method == 'POST':                  page_instance = get_object_or_404(pages, pk=page_id)     if page_id:      pages = FlatPage.objects.filter(sites__id__exact=kiosko.site.pk)      page_instance = None     kiosko = Kiosko.objects.get_current() def new_page(request, page_id=None): @user_passes_test(is_store_admin)      )         template_name='kiosquero/manage_pages.html',         pages,         request,     return object_list(          pages = FlatPage.objects.filter(sites__id__exact=kiosko.site.pk) ad     �     h       �  �  u  V  2    �  �  �  E    �  �  o  a  6    �  �  �  �  �  w  m  l  M  :    �  �  �  �  �  �  z  y  W  <    �
  �
  �
  �
  f
  4
  3
  
  �	  �	  �	  N	  9	  	  �  �  }  V  )  �  �  �  j  5    �  �  �  [  6    �  �  v  3  �  �  �  �  �  �  Z  C  4    �  �  �  ~  p  j  i  S  )  �  �  �  �  �  w  Y  8  
  �  �  �                           data = form.cleaned_data         if form.is_valid():         form = ConfigDomainForm(request.POST)     if request.method == 'POST':     form = ConfigDomainForm()     errors = []     kiosko = Kiosko.objects.get_current() def config_domain(request): @user_passes_test(has_domain)      return kiosko.plan.has_domain() and is_store_admin(user)     kiosko = Kiosko.objects.get_current() def has_domain(user):      )             }             'errors':errors,             'kiosko':kiosko,             'live_forms': live_forms,             'store_config_form': store_config,             'seller_form':seller_form,             {          extra_context=         'kiosquero/config_store.html',          request,       return direct_to_template(              errors = [_("Correct the errors below")]         else:             return HttpResponseRedirect(reverse("manage"))             cache.delete(GET_CONFIG_CACHE_KEY % {'id': kiosko.id})             store_conf.save()             store_conf.store_description = data['description_store']             store_conf = kiosko.get_config()                 return redirect('store_delete')             if data['remove_store']:             kiosko.plan = data['plan']             data = store_config.cleaned_data             # Config             request.user.message_set.create(message=_('Store configuration updated.'))             seller.save()             seller.receive_updates = data['updates']             seller.postcode = data['zipcode']             seller.city = data['city']             seller.state = data['state'].name             seller.country = data['country'].printable_name             seller.address = data['address']             seller.cuit = data['cuit']             seller.telephone = data['phone']             seller.last_name = data['sellerlastname']             seller.name = data['sellername']             data = seller_form.cleaned_data             # Seller         if seller_form.is_valid() and store_config.is_valid():          store_config = ConfigStoreForm(request.POST, kiosko=kiosko)         seller_form = SellerForm(request.POST, instance=seller)     if request.method == 'POST':      store_config = ConfigStoreForm(kiosko=kiosko)     seller_form = SellerForm(instance=seller)     live_forms = config_live(request, [GoogleSettingsForm,])     errors = []      seller = Seller.objects.from_kiosko(kiosko)     kiosko = Kiosko.objects.get_current() def config_store(request): @user_passes_test(is_store_admin)      )             }             'skins':skins             'kiosko':kiosko,             'config_form':config_form,             {          extra_context=         'kiosquero/design_store.html',          request,       return direct_to_template(          )             }                 'banner':kiosko.banner,                 'logo':kiosko.logo,             {             },             'skin':kiosko.skin,             'incountries': incountries,             'shop_name': kiosko.site.name,             {         config_form = ConfigForm(         incountries = [unicode(pk) for pk in pks]         pks = shop_config.shipping_countries.all().values_list('pk', flat=True)     if not config_form or config_form.is_valid():             request.user.message_set.create(message=_('Design of store configuration updated.'))             kiosko.save()                 kiosko.banner.delete()             if data['remove_banner']:                 kiosko.logo.delete()             if data['remove_logo']:             kiosko.site.save()             shop_config.save()                 shop_config.shipping_countries.add(country)             for country in data['incountries']: ad  0   �     ]       �  t  .  �  �  R    �  �  G    �  �  �  v  A  @  !    �  �  �  �  �  ~  x  w  U  :  1    �
  �
  
  8
  ,
  
  �	  �	  �	  R	  3	  2	  1	  	  �  �  �  k  J  %  �  �  s  n  V  E  3  �  �  �  �  {  q  k  j  H  �  �  �  �  t  ;  :  %  �  �  �  m  I    �  �  �  T  9    �  �  Y  1  �  �  �                                                                                            request.FILES,             image_form = ProductImageForm(request.POST,             rename_files(request.FILES)                                              instance=product)             attributes_form = AttributesForm(request.POST,                                    instance=product)             price_form = PriceForm(request.POST,             product.save()                 product.date_added = datetime.date.today()             if not product.pk:             # force to add the creation date             product.rubro_set = product_form.cleaned_data['rubros']             product = product_form.save()         if product_form.is_valid():         product_form = ProductForm(request.POST, instance=product_instance)     if request.method == 'POST':          product_instance = get_object_or_404(products, slug=product_slug)     if product_slug:      products = Product.objects.filter(site=kiosko.site)      product_instance = None     kiosko = Kiosko.objects.get_current()     errors = []                 special=('_tag', '../')): def new_product(request, product_slug=None, template='kiosquero/product_form.html', @user_passes_test(is_store_admin)      )         }             'state': state,             'out_of_stock':out_of_stock,             'in_stock':in_stock,         extra_context = {         template_name='kiosquero/manage_products.html',         products,         request,     return object_list(          out_of_stock = len([p for p in products if not p.in_stock])         in_stock = len([p for p in products if p.in_stock])             products = products.filter(active=active)         active = (state == 'active')     if state and state != 'all':     products = Product.objects.filter(site=kiosko.site)     kiosko = Kiosko.objects.get_current()     state = request.GET.get('state', None) def products(request): @user_passes_test(is_store_admin)                                )                               extra_context= { 'object':kiosko }                               'kiosquero/confirm_delete.html',     return direct_to_template(request,         raise Http404         # fail security test     except:             return HttpResponseRedirect("http://%s"%request.main_site)             kiosko.save()             kiosko.active = False         if request.method == 'POST' and request.POST['post'] == u"yes":         kiosko = Kiosko.objects.get_current()     try: def store_delete(request): @user_passes_test(is_store_admin)      )             }             'errors':errors,             'form': form,             {         extra_context=         'kiosquero/config_domain.html',         request,     return direct_to_template(              errors = [_("Correct the errors below")]         else:             return redirect("manage")             request.user.message_set.create(message=msg)             msg = _('Domain configuration updated.')                       to, fail_silently=False)             send_mail(subject, text, settings.DEFAULT_FROM_EMAIL,             to = [admin[1] for admin in settings.ADMINS]                                                 'plan': kiosko.plan})                                                 'domain': data['domain'],                                                 'olddomain':kiosko.site.domain,                                                 'name': kiosko.get_name(),                      'Store %(name)s has this plan %(plan)s' % {                      '%(olddomain)s to this new one %(domain)s. \n' \             text = _('Store %(name)s need to change its domain: \n'             subject = _('Domain change %(kiosko)s' % {'kiosko':kiosko}) 