b0VIM 7.3      �,-M�z �  pandres                                 acerina                                 ~pandres/projects/bixti/leonidas/apps/search/views.py                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        utf-8	 3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp	                                       P                            W       _                     @       �              	       !       �                     b                           3       y             
       3       �                           �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ad  �  \            �  �  �  �  P  /    �  �  ~  Z  '  �  �  �  ]  \  �  �  �  ~  g  f  7        �  �  q  F  "  �
  �
  �
  �
  �
  �
  g
  %
  �	  �	  �	  v	  u	  t	  N	  	  �  �  �  �  }  k  B  �  �  �  �  �  ,  +  �  �  �  N       �  �  �  k  7    �  u  t  P     �  �  �  �  �  h  @  )  �  �  �  <    �  �  �  �                # get related products           #    property_values.append(pv.value)         #for pv in product.property_value.all():         #property_values = []         #product = get_object_or_404(models.Product, pk=product_id)         product = get_object_or_404(Product, pk=product_id)         #from common.models import Product   # cometa         from product.models import Product # kioskito      if params is None:     params = cache.get(cache_key, None)     cache_key = "product_params_%s" % product_id def show_product(request, product_id, name): @cache_page(settings.PAGE_VIEW_CACHE)           context_instance=RequestContext(request))         {'latest_added':latest_added_products},     return render_to_response(tpl,           return HttpResponseRedirect(prefix+iri_to_uri('/find/%s' % query))             return HttpResponseRedirect(prefix+iri_to_uri('/find-store/%s' % query))         if search_by == 'stores':         query = query.replace('/', query_space_sep)         query = query.replace('-', query_space_sep)         query = query.replace(' ', query_space_sep)         query = slugify(query)     if query:          cache.set(latest_added_prods_key, latest_added_products, cache_time)         latest_added_products = Product.objects.all().order_by('-id')[:12]     if not latest_added_products:     latest_added_products = cache.get(latest_added_prods_key)     latest_added_prods_key = "latest_added_prods"          return HttpResponseRedirect(prefix+iri_to_uri('/property/target/%s' % targets))         targets = '-'.join(targets)      if targets:     targets = request.GET.getlist('target')          return HttpResponseRedirect(prefix+iri_to_uri('/property/material/%s' % materials))         materials = '-'.join(materials)      if materials:     materials = request.GET.getlist('material')     properties = {}      search_by = request.GET.get('search-by', '')     query = request.GET.get('search', '') def index(request, tpl="index.html", prefix=""): @cache_page(settings.PAGE_VIEW_CACHE)   come_from_store = re.compile(r'^https?://[^/]+/store/(\d)/[^/]+')  max_related = getattr(settings, "MAX_RELATED_PRODUCTS", 5) cache_time = getattr(settings, "CACHE_TIME", 60) query_space_sep = getattr(settings, 'QUERY_SPACE_SEPARATOR', '+') category_space_sep = getattr(settings, 'CATEGORY_SPACE_SEPARATOR', '-')  log = get_logger('bixti.search.views')  from logger import get_logger   from heladera.models import Kiosko, Rubro from product.models import Category from common.models import Country, Partner from common import models from product.models import Product, AttributeOption, ProductAttribute from perseidas.updater.single_update import update_product    from livesettings.models import Setting from livesettings import ConfigurationSettings          currencysymbol from leonidas.apps.search.templatetags.search_extras import escape_category,\ from leonidas.apps.utils.views import get_pag  @c  @cache_page_with_prefix(60*15, lambda request: md5_constructor(str(request.GET)).hexdigest()) from django.utils.hashcompat import md5_constructor from view_cache_utils import cache_page_with_prefix from django.views.decorators.cache import cache_page from django.utils.encoding import iri_to_uri from django.utils.translation import ugettext as _ from django.utils import simplejson from django.core.cache import cache from django.shortcuts import get_object_or_404 from django.template.defaultfilters import slugify from django.template import RequestContext from django.forms import widgets from django.template.defaultfilters import urlencode from django.http import HttpResponseRedirect, Http404, HttpResponse from django.conf import settings import re import math ad  A  m            �  �  n  m  l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  context_instance=RequestContext(request))     return render_to_response('specials.html', {}, def specials(request): ad    �     P       �  �  W  	  �  �  �  t  L  J  I    �  �  �  _  5  4      �  �  �  b  1  �  �  �  �  �  �  Z  0  �
  �
  �
  �
  �
  
  #
  "
  �	  �	  �	  i	  h	  6	  �  �  �  >  =  /    �  �  t  R  �  �  �  �  ]  +  *  )    �  �  }  f  /  �  �  y  [  *  �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             # get related products           #    property_values.append(pv.value)         #for pv in product.property_value.all():         #property_values = []         #product = get_object_or_404(models.Product, pk=product_id)         product = get_object_or_404(Product, pk=product_id)         #from common.models import Product   # cometa         from product.models import Product # kioskito      if params is None:     params = cache.get(cache_key, None)     cache_key = "product_params_%s" % product_id def show_product(request, product_id, name): @cache_page(settings.PAGE_VIEW_CACHE)           context_instance=RequestContext(request))         {'latest_added':latest_added_products},     return render_to_response(tpl,           return HttpResponseRedirect(prefix+iri_to_uri('/find/%s' % query))             return HttpResponseRedirect(prefix+iri_to_uri('/find-store/%s' % query))         if search_by == 'stores':         query = query.replace('/', query_space_sep)         query = query.replace('-', query_space_sep)         query = query.replace(' ', query_space_sep)         query = slugify(query)     if query:          cache.set(latest_added_prods_key, latest_added_products, cache_time)         latest_added_products = Product.objects.all().order_by('-id')[:12]     if not latest_added_products:     latest_added_products = cache.get(latest_added_prods_key)     latest_added_prods_key = "latest_added_prods"          return HttpResponseRedirect(prefix+iri_to_uri('/property/target/%s' % targets))         targets = '-'.join(targets)      if targets:     targets = request.GET.getlist('target')          return HttpResponseRedirect(prefix+iri_to_uri('/property/material/%s' % materials))         materials = '-'.join(materials)      if materials:     materials = request.GET.getlist('material')     properties = {}      search_by = request.GET.get('search-by', '')     query = request.GET.get('search', '') def index(request, tpl="index.html", prefix=""): @cache_page(settings.PAGE_VIEW_CACHE)   come_from_store = re.compile(r'^https?://[^/]+/store/(\d)/[^/]+')  max_related = getattr(settings, "MAX_RELATED_PRODUCTS", 5) cache_time = getattr(settings, "CACHE_TIME", 60) query_space_sep = getattr(settings, 'QUERY_SPACE_SEPARATOR', '+') category_space_sep = getattr(settings, 'CATEGORY_SPACE_SEPARATOR', '-')  log = get_logger('bixti.search.views')  from logger import get_logger   from heladera.models import Kiosko, Rubro from product.models import Category from common.models import Country, Partner from common import models from product.models import Product, AttributeOption, ProductAttribute from perseidas.updater.single_update import update_product    from livesettings.models import Setting from livesettings import ConfigurationSettings          currencysymbol from leonidas.apps.search.templatetags.search_extras import escape_category,\ from leonidas.apps.utils.views import get_page, get_letter_list, find_setting from leonidas.indexservice.client import IndexProduct, OR_OPERATOR from leonidas.apps.paginator import CustomPaginator from leonidas.shortcuts import render_to_response ad  �  �     3       �  �  �  1    �  �  �  �  x  <  �  �  �  �    ~  u  H      �  �  z  e  d  H  ,    �  �  {  A  )  �
  �
  �
  u
  Y
  7
  
  
  �	  �	  �	  ~	  K	  	  	  	  �  �  i  m  Q    �  �  n  m  ^  U  #    �  �  �  �  �  �  Z    �  �  �  �    =  �  �  �  �  q  U    �  �  �  �  b  [  (  �  �  �  �  �  U  T  8    �  �                                      'category_list.html',(), filter_by={'parent': None})     return get_letter_list(request, Rubro, def category_list(request):                   'brands_list.html', ('id', 'name', 'logo'))     return get_letter_list(request, models.Brand, def brands_list(request):                                 context_instance=RequestContext(request))     return render_to_response(tpl, initial_params,     })         'search_by_store': True,         'partner_id': request.partner_id,         'raw_query': raw_query or '',         'get': get and get + "&",         'query': search_text or '',         'sort_widget': sort_widget.render('sort', sort_by),         'time': index.time,         'results': results,     initial_params.update({                                            ('>price', _('Mayor Precio'))])                                           ('<price', _('Menor Precio')),     sort_widget = widgets.Select(choices=[('', _('Relevancia')),                         for x, y in request.GET.iteritems() if x != 'p'))     get = '&'.join(("%s=%s" % (x, y ) #and y[0])       results = paginator.page(page)     paginator = CustomPaginator(index, slimit, psize=limit)     index = IndexProduct(search_str=search_text, store_name=True)          page = 1     except ValueError:         page = int(request.GET.get('p', 1))     try:         limit = 1     except ValueError:         limit = int(request.GET.get('l', slimit))     try:     slimit = 6                      else ('score', False)     tsort_by = (sort_by[1:], sort_by.startswith('>')) if sort_by \     sort_by = request.GET.get('sort', '')     search_text = search_text and search_text.replace(query_space_sep, ' ')     raw_query = search_t@cache_page_with_prefix(settings.PAGE_@@cache_page_with_prefix(settings.PAGE_VIEW_CACHE, lambda request: md5_constructor(str(request.GET)).hexdigest())                                 context_instance=RequestContext(request))     return render_to_response(tpl, initial_params,     })         'partner_id': request.partner_id,         'raw_query': raw_query or '',         'product_materials': product_materials,         'zones': zones,         'fzones': fzones,         'filterscat': filterscat,         'filters': filters,         'get': get and get + "&",         'query': search_text or '',         'price_range': {'from': price_from, 'to': price_to},         'in_brands': '', #search_text in brands,         'rubro': rubro,         'category': escape_category(category), #category,         'categories': categories,         'top_level': 1, # if lvl is None else lvl + 2,         'sort_widget': sort_widget.render('sort', sort_by),         'time': index.time,         'results': results,     initial_params.update({          rubro = None     except Exception, e:             cache.set(cache_key, rubro, cache_time)             rubro = Rubro.objects.get(name__icontains=category)         if not rubro:         rubro = cache.get(cache_key, None)         cache_key = "rubro_%s" % (category,)     try:              product_materials.append(attrib.value)         if attrib.name == 'material':     for attrib in product_attributes:          cache.set(cache_key, product_attributes, cache_time)         product_attributes = ProductAttribute.objects.all()     if not product_attributes:     product_attributes = cache.get(cache_key, None)     cache_key = "product_attributes"      product_materials = []     #    cache.set("brands", brands)     #    brands = [b["search_term"].replace(query_space_sep,' ') for b in brands]     #    brands = models.Brand.objects.values("search_term")     #if brands is None:     #brands = cache.get("brands", None) ad     �     b       �  �  d  "  �  �  �  �  �  i  `  .      �  �  �  �  �  �  ]  6      �  �  �  d  /  �  �  �  J      �
  �
  �
  S
  "
  �	  �	  �	  �	  <	  	  �  �  �  {  K    �  q  ,  �  �  �  �  s  H  .  -      �  �  �  e  V  U  D  3    �  �  �  �  a  :  /  *    �  �  �  [  P  O    �  z  y  G  �  �  �  �  �                    filterscat = filter(lambda x: x.get("filter", "")=="category", filters)                        for x, y in request.GET.iteritems() if x != 'p'))     get = '&'.join(("%s=%s" % (x, y ) #and y[0])                                             ('>price', _('Mayor Precio'))])                                           ('<price', _('Menor Precio')),     sort_widget = widgets.Select(choices=[('', _('Relevancia')),           })                            _('a') + " $%d " % price_to,             'description': _('De') + " $%d " % price_from + \             'filter': 'price_from,price_to',         filters.append({     if price_from:              })             'description': cat_filter,             'filter': 'category',          filters.append({         #        cat_filter = cat         #    if escape_category(cat) == category:         #for lv, cat in categories:         cat_filter = category     if category:     filters = []              })                 'description': "%s"%state['name'],                 'filter': 'state-%s'%state['clean_name'],              fzones.append({         for state in vstates:     if vstates:     fzones = []      #categories.reverse()     #                     actual=category)     #lvl = get_categories(index.categories.items(), res=categories,      categories = []      results = paginator.page(page)     paginator = CustomPaginator(index, slimit, psize=limit)                          properties=properties, category_name=rubro)                          sort_by=tsort_by, store=store, states=states,                           price_from=conv_price_from, price_to=conv_price_to,     index = IndexProduct(search_str=search_text, category=category,      #    not initial_params and not properties:     #if not search_text and not store and not rubro and \      else: conv_price_to = None     if price_to>=0: conv_price_to = price_to*float(conversion_rate)+1     else: conv_price_from = None     if price_from>=0: conv_price_from = price_from*float(conversion_rate)                    (conversion_rate, symbol), cache_time)         cache.set("currency_%s" % request.country_id,             "default_currency__symbol",)[0]             "default_currency__conversion_rate",         conversion_rate, symbol = country.values_list(              cache.set(cache_key, country, cache_time)             country = Country.objects.filter(pk=request.country_id)         if not country:         country = cache.get(cache_key, None)         cache_key = "country_%s" % (request.country_id,)     if not conversion_rate or not symbol:                                         (None, None))     conversion_rate, symbol = cache.get("currency_%s" % request.country_id,     # Convert prices from default country's currency     if price_to and not price_from: price_from = 0         price_to = None     except (TypeError, ValueError), e:         price_to = int(request.GET.get('price_to')) #or None     try:         price_from = None     except (TypeError, ValueError), e:         price_from = int(request.GET.get('price_from')) #or None     try:          page = 1     except ValueError:         page = int(request.GET.get('p', 1))     try:         limit = 1     except ValueError:         limit = int(request.GET.get('l', slimit))     try:     slimit = settings.DEFAULT_PAGINATE_BY      #        states = None     #        vstates = []     #    except:     #        states = " ".join([str(state['id']) for state in vstates])     #        vstates = pstates.values('name', 'clean_name', 'id')     #            pstates = pstates.exclude(clean_name=state)     #        for state in excluded_states:     #        zones = pstates = partner.states.all() ad  �  �     @       �  �  �  r  q  ^  >    �  �  �  q  A  #  �  �  �  �  �  R  H      �  �  �  g  4  �  �  �  g    �
  �
  
  ~
  C
  �	  �	  �	  �	  �	  [	  Z	  	  �  �  �  g  [  A    �  �  l  k  �  �  �  e  d  c  �  �  �  �  �  �  �  f  ?  >    �  �  Q  &  %    �  �  }  :    �  �  �  �  �  �  ^  ,    
  �  �  �                                #        partner = Partner.objects.get(id=request.partner_id)     #    try:     #if not store:     zones = []     #excluded_states = excluded_states.split('-')     #excluded_states = request.GET.get('exclude', "")     states = None     vstates = []     # filter by states using partner                          # else ('date_added', True)                    else ('score', False)     tsort_by = (sort_by[1:], sort_by.startswith('>')) if sort_by \     sort_by = request.GET.get('sort', '')     search_text = search_text and search_text.replace(query_space_sep, ' ')     raw_query = search_text     #    return match      #        res.append((level, category))     #        match = actualm or (level if normcat == actual else None)     #        normcat = escape_category(category)     #        actualm = get_categories(sub.items(), res, level + 1, actual)     #    for category, sub in categories:      #    categories.sort(reverse=True)     #    # Sort level alphabetically      #        return     #    if not categories:     #def get_cat@cache_page_with_prefix(settings.PAGE_@cache_page_with_prefix(settings.PAGE_VIEW_CACHE, lambda request: md5_constructor(str(request.GET)).hexdigest())       return search(request, '', '', properties={propty:values})     values = values.replace('-', ' ') def search_properties(request, propty, values): @cache_page_with_prefix(settings.PAGE_VIEW_CACHE, lambda request: md5_constructor(str(request.GET)).hexdigest())                          mimetype='application/javascript')     return HttpResponse(simplejson.dumps(price),               'currency': currencysymbol(dproduct['store__country']),}     price = {'price': finalprice,         finalprice = None     except:         finalprice = str(uproduct['properties'][56])     try:     uproduct = update_product(dproduct)                 'store': product.store.id, 'url': product.url}     dproduct = {'id': product.id, 'store__country': product.store.country.id,      cache.delete("cluster_%s"%product.cluster.id)     product = get_object_or_404(models.Product, pk=product_id) def ajax_product_price(request, product_id):                                 context_instance=RequestContext(request))     return render_to_response('show_product.html', params,      #        return HttpResponseRedirect(url)     #           params['partner_id'])     #           product.store_id, params['cluster'].type_id or "",     #           urlencode(product.url), slugify(product.store.name), product.id,     #        url = "/redirect/?url=%s&sname=%s&pid=%s&stid=%s&tid=%s&paid=%s"%(     #        product = product[0]     #    if len(product) == 1:     #                    if p.store_id == int(store_id[0])]     #    product = [p for p in params['products']      #if len(store_id) == 1:     #store_id = come_from_store.findall(referer)     #referer = request.META.get('HTTP_REFERER', '')     # if comming from store redirect to store          cache.set(cache_key, params, cache_time)         }             'partner_id': request.partner_id,              # Tracking             'tags': tags,             'targets': targets,             'materials': materials,             'total_products':total_products,             'rubros': rubros,             'prod_categories': prod_categories,             'categories': categories,             'shippings': shippings,             'payments': payments,             'featured_products':featured_products,             'product_kiosko': product_kiosko,             'product': product,         params = {              log.error('Can not get shippings from product %s, error: %s'%(product, e))         except Exception, e:                      pass ad     �     W       �  v  u  8    �  �  �  o  @        �  �  �  u  F    �  �  �  �  �  O  2      �  �  �  �  v  4  �
  �
  �
  O
  N
  *
  
  
  �	  }	  N	  &	  		  �  �  �  �  ;    �  �  �  O  '  �  �  �  Y    �  �  �  ,  +  �  �  �  n  D  �  �  �  �  /  �  �  �  �  �  D  �  �  �  �                               except:                     shippings[method] = ' - $'.join([shippings[method], m_rate])                                        site=product_kiosko.site, default=False).value                     m_rate = find_setting('SHIPPING', '%s_RATE'%(method_keyword,),                  try:                      pass                 except:                     shippings[method] = ' - '.join([shippings[method], m_days])                                            site=product_kiosko.site, default=False).value                     m_days = find_setting('SHIPPING', '%s_DAYS'%(method_keyword,),                  try:                          _(u"Per unit shipping fee: {label}".format(label=label))                     shippings[method] = \                 else:                         _(u"General shipping fee: {label}".format(label=label))                     shippings[method] = \                 if method_keyword == 'FLAT':                  label = find_setting('SHIPPING', method, site=product_kiosko.site).value                 method = method_keyword+'_SERVICE'                 method_keyword = shipping.split('.')[-1].upper()             for shipping in modules:             #modules = unicode(modules).replace('\'', '"')             #log.debug("modules: %s - type: %s",modules, type(modules))                  modules = simplejson.loads(modules)                 modules = unicode(modules).replace('\'', '"').replace("[u", "[")                 modules = modules.value             if modules and type(modules) != list:                                                 site=product_kiosko.site, default=True)             modules = find_setting('SHIPPING', 'MODULES',              # needs heavy refactoring.             # this section, and maybe the previous too, together with find_setting         try:         shippings = {}              log.error('Can not get payments from product %s, error: %s'%(product, e))         except Exception, e:             # get Shipping from product                 payments[payment.slug] = label                 label = find_setting(payment.slug, 'LABEL', site=site_id).value             for payment in product_kiosko.payments.all():         try:         payments = {}         # get Payments from product              cache.set(prod_tot_key, str(total_products), cache_time)             total_products = Product.objects.filter(site=site_id).count()         if not total_products:         total_products = cache.get(prod_tot_key, None)         prod_tot_key = "total_products_site_idex_%s" % (site_id,)                          featured=True)[:6]         featured_products = Product.objects.filter(site=site_id, \          site_id = product_kiosko.site_id              product_kiosko = None         except Exception, e:             product_kiosko = product.site.kiosko_set.all()[0]         try:                  tags.append(attrib.value)             elif attrib.name == u'tags':                 targets.append(attrib.value)             elif attrib.name == u'target':                 materials.append(attrib.value)             if attrib.name == u'material':         for attrib in product.productattribute_set.all():         tags = []         targets = []         materials = []          #    rubros.append(rubro.name)         #for rubro in product.rubro_set.all():         rubros = []          prod_categories = product.category.all()         categories = Category.objects.filter(site=product.get_kiosko().site)         #            if idx.cluster_id != cluster_id]         #related = [idx for idx in index[:max_related + 1] \          #                     default_operator=OR_OPERATOR)         #index = IndexProduct(search_str=product.name, get_categories=False,  ad  �
  2     !       �  r  4        �  �  �  �  A    �  �  �  �  k    �  �  �  Z  U  T  /      �  �  �  �  t  2  
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                #        partner = Partner.objects.g    #        partner = Partner.objects.get(id=request.partner_id)     #    try:     #if not store:     zones = []     #excluded_states = excluded_states.split('-')     #excluded_states = request.GET.get('exclude', "")     states = None     vstates = []     # filter by states using partner                          # else ('date_added', True)                    else ('score', False)     tsort_by = (sort_by[1:], sort_by.startswith('>')) if sort_by \     sort_by = request.GET.get('sort', '')     search_text = search_text and search_text.replace(query_space_sep, ' ')     raw_query = search_text     #    return match      #        res.append((level, category))     #        match = actualm or (level if normcat == actual else None)     #        normcat = escape_category(category)     #        actualm = get_categories(sub.items(), res, level + 1, actual)     #    for category, sub in categories:      #    categories.sort(reverse=True)     #    # Sort level alphabetically      #        return     #    if not categories:     #def get_categories(categories, res, level=0, actual=''):              initial_params={}, properties={}, tpl='search_results.html'): def search(request, category, search_text, store=None, rubro=None, ad    �     3       �  �  w  +    �  �  �  �  {  I  2       �  �  �  �  �  D  !     �  �  �  c    �  �  �  �  {  ?    �
  �
  �
  �
  �
  N
  
  
  
  �	  �	  {	  z	  ^	  3	  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            'category_list.html',(), filter_by={'parent': None})     return get_letter_list(request, Rubro, def category_list(request):                   'brands_list.html', ('id', 'name', 'logo'))     return get_letter_list(request, models.Brand, def brands_list(request):                                 context_instance=RequestContext(request))     return render_to_response(tpl, initial_params,     })         'search_by_store': True,         'partner_id': request.partner_id,         'raw_query': raw_query or '',         'get': get and get + "&",         'query': search_text or '',         'sort_widget': sort_widget.render('sort', sort_by),         'time': index.time,         'results': results,     initial_params.update({                                            ('>price', _('Mayor Precio'))])                                           ('<price', _('Menor Precio')),     sort_widget = widgets.Select(choices=[('', _('Relevancia')),                         for x, y in request.GET.iteritems() if x != 'p'))     get = '&'.join(("%s=%s" % (x, y ) #and y[0])       results = paginator.page(page)     paginator = CustomPaginator(index, slimit, psize=limit)     index = IndexProduct(search_str=search_text, store_name=True)          page = 1     except ValueError:         page = int(request.GET.get('p', 1))     try:         limit = 1     except ValueError:         limit = int(request.GET.get('l', slimit))     try:     slimit = 6                      else ('score', False)     tsort_by = (sort_by[1:], sort_by.startswith('>')) if sort_by \     sort_by = request.GET.get('sort', '')     search_text = search_text and search_text.replace(query_space_sep, ' ')     raw_query = search_text                  tpl='search_results_store.html'): def search_store(request, search_text, initial_params={}, 