b0VIM 7.3      q�0Mz  -  pandres                                 acerina                                 ~pandres/projects/bixti/leonidas/urls.py                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          	 3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           ^                     ��������K       _                     	       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ad     �     ^       �  �  |  G  F    �  �  �  �  �  �  �  r  V  5    �  �  �  �  �  t  =  �  �  �  �  �  ^  0  �  �  q  @  ?    �
  �
  �
  4
  �	  p	  o	  =	  �  �  �    9    �  �  0  �  �  6  4  3  2    �  �  �  �  �  d  ^  ]  \  M    �  �  �  h  5  3    �  Y  W  V  :  �  �  �  `  _  3    �  �  �  �                                       {'template': 'store_redirect.html'}),     ('^redirect/$', direct_to_template,  #        {'template': 'categories.html'}), #    ('^categories/$', direct_to_template,           {'template': 'registration/registration_done.html'}),     ('^user/register/done/$', direct_to_template,          {'login_url': LOGIN_URL}),     ('^user/logout/$', 'django.contrib.auth.views.logout_then_login', urlpatterns += patterns('',  )     ('^user/register/$','bixti_registration.views.bixti_register', {}, 'register'),     ('^user/login_then_signup/$','bixti_registration.views.login_then_signup', {}, 'login_then_signup'), urlpatterns += patterns('',  )     ('^user/crop/$', 'crop'), # move to accounts ?     ('^user/rate/$', 'rate'), # move to accounts ?     ('^user/register/confirm/$', 'activate'),     ('^user/profile/$','show_profile'),   #  ('^user/login/$', 'show_login'),  urlpatterns += patterns('leonidas.apps.users.views', # User actions       )         (r'^500.html/', 'leonidas.apps.utils.views.server_error'),     urlpatterns += patterns('', if settings.DEBUG:  )     (r'^fbyopeo/', include('leonidas.apps.fbapp.urls')), urlpatterns += patterns('',   )     #(r'^shop/contact/', 'leonidas.apps.contacts.views.shop_contact', {}, 'shop_contact'),     #    {'template':'contacts/contact_thanks.html'},'shop_contact_thanks'),     #(r'^contacto-tienda/grx/$','django.views.generic.simple.direct_to_template',     (r'^contacto-tienda/', 'leonidas.apps.contacts.views.shop_contact', {}, 'shop_contact'),     url(r'^media/skins/style.css', 'kiosquero.views.skin_css', name='skin_css'),     (r'^cart/', include('global_cart.urls')),     (r'^captcha/', include('captcha.urls')),         {'document_root': settings.MEDIA_ROOT, 'show_indexes':True}),     (r'^media/(?P<path>.*)$', 'django.views.static.serve',      (r'^admin/', include(admin.site.urls)),      url(r'^user-login/$', 'bixti_registration.views.shop_login', name='user_login'),     (r'^accounts/', include('multicuenta.urls')),      url(r'^manage/section/(?P<category_slug>[^/]+)/$','kiosquero.views.new_category', name='edit_category'),     url(r'^manage/section/add/$','kiosquero.views.new_category', name='new_category'),     url(r'^manage/section/$', 'kiosquero.views.category', name='categories'),      url(r'^manage/credit/$', 'multicuenta.views.user_account', name='multicuenta_user_account'),     (r'^manage/', include('featured.urls')),     (r'^manage/', include('kiosquero.urls')),      (r'^mostrador/', include('mostrador.urls')),     url(r'^shop/logout/$', 'mostrador.views.shop_logout', name='shop_logout'),         name='redirect_to_account'),     url(r'^redirect-to-account/$', 'mostrador.views.redirect_to_account',      (r'^product/', 'mostrador.views.signup'),     (r'^signup/', 'mostrador.views.signup'), urlpatterns += patterns('',  )     (r'^blank_base/$', 'direct_to_template', {'template': 'base.html'}),     (r'^blank/$', 'direct_to_template', {'template': 'base_blank.html'}), urlpatterns += patterns('django.views.generic.simple', #if settings.DEBUG:  handler404 = 'leonidas.apps.utils.views.not_found' handler500 = 'leonidas.apps.utils.views.server_error'  SUCCESS_REGISTER_URL = PROFILE_URL PROFILE_URL = '/user/profile/' FORGOT_PWD_URL = '/user/forgot/' #LOGIN_URL = '/user/login/' RATE_URL = '/user/rate/' ACTIVATION_URL = '/user/register/confirm/' # useful urls  admin.autodiscover() from django.contrib import admin  from settings import LOGIN_URL from satchmo_store.urls import urlpatterns  from django.views.decorators.cache import cache_page from django.views.generic.simple import direct_to_template from django.conf.urls.defaults import * from django.conf import settings ad  j  �     	       �  �  �  �  f  /  �  �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ) #        ('^review/create/$', 'leonidas.apps.users.views.create_review'),             {'document_root': settings.MEDIA_ROOT}),         (r'^media/(.*)$', 'django.views.static.serve',     urlpatterns += patterns('', if settings.DEBUG:  )     url('^rubros/(?P<rubro>[\w-]+)/$', 'search', {'search_text':'', 'category':''}, name='search'), 